`include "uvm_pkg.sv"
package adder_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "sequence_item.sv"
    `include "sequence.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent_config.sv"
    `include "agent.sv"
    `include "scoreboard.sv"
    `include "env_config.sv"
    `include "environment.sv"
    `include "test.sv"

endpackage : adder_pkg