`define DATA_WIDTH 16
`define ADDR_WIDTH 8
`define DEPTH 256
`define RESET_VALUE 16'h5678