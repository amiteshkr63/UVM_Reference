`include "uvm_pkg.sv"
package memory_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "memory_seq_item.sv"
    `include "memory_sequence.sv"
    `include "memory_driver.sv"
    `include "active_memory_monitor.sv"
    `include "passive_memory_monitor.sv"
    `include "active_memory_agent.sv"
    `include "passive_memory_agent.sv"
    `include "memory_scoreboard.sv"
    `include "memory_environment.sv"
    `include "memory_test.sv"
endpackage : memory_pkg